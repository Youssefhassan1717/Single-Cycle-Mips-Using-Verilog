`timescale 1ns / 1ps

module InstructionMemory(
    input CLK,
    input [31:0] Address,
    output reg [31:0] Instr
    );
    
reg [31:0] ROM [0:2147483648];

initial 
    begin
    
        //Test case 0
        ROM[0] = 32'b00100000000100000000000000000100; //ADDI $s0, $zero, 4
        ROM[1] = 32'b00100000000100010000000000000011; //ADDI $s1, $zero, 3
        ROM[2] = 32'b00000010000100011001000000100101; //OR $s2, $s0, $s1
        
        //Test case 1
        ROM[4] = 32'b00100000000100000000000000000001; //ADDI $s0, $zero, 1
        ROM[5] = 32'b00100000000100010000000000000011; //ADDI $s1, $zero, 3
        ROM[6] = 32'b00000010001100001001000000100100; //AND $s2, $s1, $s0
        
        //Test case 2
        ROM[8] = 32'b00100000000100001111111111111111; //ADDI $s0, $zero, 65535
        ROM[9] = 32'b00100000000100010000000000000001; //ADDI $s1, $zero, 1
        ROM[10] = 32'b00000010001100001001000000100000; //ADD $s2, $s1, $s0
        
        //Test case 3
        ROM[12] = 32'b00100000000100000000000000001000; //ADDI $s0, $zero, 8
        ROM[13] = 32'b00100000000100010000000000000001; //ADDI $s1, $zero, 1
        ROM[14] = 32'b00000010000100011001000000100010; //SUB $s2, $s0, $s1
        
        //Test case 4
        ROM[16] = 32'b00100000000100000000000000000101; //ADDI $s0, $zero, 5
        ROM[17] = 32'b00100000000100010000000000000100; //ADDI $s1, $zero, 4
        ROM[18] = 32'b00000010001100001001000000100000; //ADD $s2, $s1, $s0
        
        //Test case 5
        ROM[20] = 32'b00100000000100000000000001100100; //ADDI $s0, $zero, 100
        ROM[21] = 32'b00100000000100010000000111110100; //ADDI $s1, $zero, 500
        ROM[22] = 32'b00000010000100011001000000100010; //SUB $s2, $s0, $s1
    
   end
    
always @(posedge CLK)
    begin
        Instr <= ROM[Address];
    end
    
endmodule
